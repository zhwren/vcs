/*******************************************************************************
**                                  _ooOoo_                                   **
**                                 o8888888o                                  **
**                                 88" . "88                                  **
**                                 (| -_- |)                                  **
**                                  O\ = /O                                   **
**                              ____/`---'\____                               **
**                            .   ' \\| |// `.                                **
**                             / \\||| : |||// \                              **
**                           / _||||| -:- |||||- \                            **
**                             | | \\\ - /// | |                              **
**                           | \_| ''\---/'' | |                              **
**                            \ .-\__ `-` ___/-. /                            **
**                         ___`. .' /--.--\ `. . __                           **
**                      ."" '< `.____<|>_/___.' >'"".                         **
**                     | | : `- \`.;` _ /`;.`/ - ` : | |                      **
**                       \ \ `-. \_ __\ /__ _/ .-` / /                        **
**               ======`-.____`-.___\_____/___.-`____.-'======                **
**                                  `=---='                                   **
**                                                                            **
**               .............................................                **
**                      Buddha bless me, No bug forever                       **
**                                                                            **
********************************************************************************
** Author           :     ZhuHaiWen                                           **
** Email            :     zhuhw@ihep.ac.cn/zhwren0211@whu.edu.cn              **
** Last modified    :     2022-07-02 20:18:00                                 **
** Filename         :     test.sv
** Phone Number     :     18625272373                                         **
** Discription      :                                                         **
*******************************************************************************/
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "env.sv"

module test;
    initial begin
        run_test("env");
    end
endmodule
